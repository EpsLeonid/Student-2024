`ifndef PARAMS_v_6
`define PARAMS_v_6

package package_settings_v_6;

	parameter int l_v_6 = 6;
	parameter int k_v_6 = 13;
	parameter int m1_v_6 = 16;
	parameter int m2_v_6 = 1;

endpackage

`endif 