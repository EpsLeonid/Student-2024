`ifndef PARAMS_SVH
`define PARAMS_SVH

parameter WIDTH_A = 8;     
parameter WIDTH_B = 8;     
parameter WIDTH_C = 8;     
parameter WIDTH_OUT = 16;  

`endif
