`ifndef PARAMS_V_1
`define PARAMS_v_1
package package_settings_v_1;
    parameter int k_v_1 = 8;    
    parameter int l_v_1 = 5;    
    parameter int M_v_1 = 16;   
endpackage
`endif