`ifndef PARAMS_V_2
`define PARAMS_V_2
package package_settings_v_2;
	parameter int k_v_2 = 5;
	parameter int l_v_2 = 5;
	parameter int M_v_2 = 16;
endpackage
`endif