`ifndef PARAMS_V5
`define PARAMS_V5

package package_settings_v_5;

	parameter int k_v_5 = 6;
	parameter int l_v_5 = 6;
	parameter int M_v_5 = 16;

endpackage

`endif