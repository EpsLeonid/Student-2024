`ifndef PARAMETER
`define PARAMETER

parameter int WIDTH = 8;
parameter int OUT_WIDTH = 2*WIDTH;

`endif