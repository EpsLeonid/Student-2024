`ifndef PARAMS_SV
`define PARAMS_SV

package package_settings_v_5;
//-----------------------------------------------------------------------------
// Parameter Declaration(s)
//-----------------------------------------------------------------------------
	parameter int k_v_5 = 6;
	parameter int l_v_5 = 6;
	parameter int M_v_5 = 16;
//-----------------------------------------------------------------------------
endpackage

`endif // PARAMS_SV