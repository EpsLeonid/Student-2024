`ifndef PARAMS_SV
`define PARAMS_SV

package params;
    parameter int DATA_WIDTH = 8; // ������ ������ A, B, C
    parameter int DATA_OUT_WIDTH = DATA_WIDTH * 2; // ������ �������� ������
endpackage

`endif // PARAMS_SV
