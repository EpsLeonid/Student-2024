`ifndef SETTINGS_v3
`define SETTINGS_v3

package package_settings_v_3;

	parameter int l_v_3 = 5;
	parameter int k_v_3 = 11;
	parameter int m1_v_3 = 16;
	parameter int m2_v_3 = 1;

endpackage

`endif 