`ifndef PARAMS_SV
`define PARAMS_SV

package package_settings_v_4;
//-----------------------------------------------------------------------------
// Parameter Declaration(s)
//-----------------------------------------------------------------------------
	parameter int k_v_4 = 9;
	parameter int l_v_4 = 5;
	parameter int M_v_4 = 16;
//-----------------------------------------------------------------------------
endpackage

`endif // PARAMS_SV